/*
*	cayde top module
*/

module cayde  ( input logic PC,
		input logic 
